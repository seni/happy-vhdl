To generate VHDL code from a grammar use the -h option.

There are two examples in examples/vhdl.
